`timescale 1ns / 1ps
//The mod flag is encoded as:
//
//Table 5.1.3: mod flag encoding
//mod bits 	description 	range of values
//	0-1 		mod.mem flag 		0-3
//	2-3 		mod.shift flag 	0-3
//	4-7 		mod.cond flag 		0-15
module instr_mod(
    );


endmodule
